package CONSTANTS is
	constant NumBit : integer := 16;	
	
end package CONSTANTS;
